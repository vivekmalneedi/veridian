module test ([5:0] clk);
endmodule


module test (logic clk);
endmodule
