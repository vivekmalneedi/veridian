module test;
  logic [1:0] abc;

  assign abc[2] = 1'b0;
endmodule
