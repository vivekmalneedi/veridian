interface simple_bus;
    logic clk;
endinterface

module test2;
    simple_bus b ();
endmodule
