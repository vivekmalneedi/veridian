module test;
    simple_bus bus ();
endmodule
