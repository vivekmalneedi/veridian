module test;
    logic abc;
    logic abcd;

  a
endmodule

