`timescale 1ns/1ps
`include "simple_bus.svh"

module test;
    simple_bus bus ();
endmodule
